configuration player_two_rgb_rom_rtl_cfg of player_two_rgb_rom is
   for rtl
   end for;
end player_two_rgb_rom_rtl_cfg;
