configuration player_pixel_mux_rtl_cfg of player_pixel_mux is
   for rtl
   end for;
end player_pixel_mux_rtl_cfg;
