configuration rom_controller_gpu_rtl_cfg of rom_controller_gpu is
   for rtl
   end for;
end rom_controller_gpu_rtl_cfg;
