configuration map_collision_checker_behavioural_cfg of map_collision_checker is
   for behavioural
   end for;
end map_collision_checker_behavioural_cfg;
