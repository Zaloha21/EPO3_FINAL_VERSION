configuration datalatchcontrol_behaviour_cfg of datalatchcontrol is
   for behaviour
   end for;
end datalatchcontrol_behaviour_cfg;
