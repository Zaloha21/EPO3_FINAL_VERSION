configuration sprite_rom_map_rtl_cfg of sprite_rom_map is
   for rtl
   end for;
end sprite_rom_map_rtl_cfg;
