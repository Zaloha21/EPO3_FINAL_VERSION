configuration movecontroller_behaviour_cfg of movecontroller is
   for behaviour
   end for;
end movecontroller_behaviour_cfg;
