library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

architecture rtl of map_rom is

    type rom_type is array (0 to 29) of std_logic_vector(39 downto 0);

	constant rom : rom_type := (
		0 => "1111111111111111111111111111111111111111",
		1 => "1000000000000000000000000000000000000001",
		2 => "1000000000000000000000000000000000000001",
		3 => "1000000000000000000000000000000000000001",
		4 => "1111111111111111111111111111111111111111",
		5 => "1000000000000000000000000000000000000001",
		6 => "1000000000000000000000000000000000000001",
		7 => "1000000000000000000000000000000000000001",
		8 => "1000000000000000000000000000000000000001",
		9 => "1110000000011111000000001111100000000111",
		10 => "1000000000010000000000000000100000000001",
		11 => "1000000111110000000000000000111110000001",
		12 => "1000000000000000000000000000000000000001",
		13 => "1000000000000000110000110000000000000001",
		14 => "1000000000000000000000000000000000000001",
		15 => "1000000000000000000000000000000000000001",
		16 => "1000111000000000000000000000000001110001",
		17 => "1000000111000000000000000000001110000001",
		18 => "1000000000000000000110000000000000000001",
		19 => "1000000000000000111001110000000000000001",
		20 => "1000000000000000000000000000000000000001",
		21 => "1110000000000000000000000000000000000111",
		22 => "1000000000010000000000000000100000000001",
		23 => "1000000000010000000000000000100000000001",
		24 => "1000000111111100000000000011111110000001",
		25 => "1000000000000000000000000000000000000001",
		26 => "1000000000000000000000000000000000000001",
		27 => "1000000000000000000110000000000000000001",
		28 => "1000000000000000011111100000000000000001",
		29 => "1111111111111111111111111111111111111111");

begin

    -- Synchronized Output
    process (clk) is
    begin
        if rising_edge(clk) then 
            if reset = '1' then
                row_of_blocks <= (others => '0');
            else 
                row_of_blocks <= rom (to_integer(unsigned(address)));
            end if;
        end if;
    end process;

end architecture rtl;