configuration player_one_sprite_rom_rtl_cfg of player_one_sprite_rom is
   for rtl
   end for;
end player_one_sprite_rom_rtl_cfg;
