configuration dataclockcontrol_behaviour_cfg of dataclockcontrol is
   for behaviour
   end for;
end dataclockcontrol_behaviour_cfg;
