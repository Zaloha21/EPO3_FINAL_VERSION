configuration bullet_controller_one_rtl_cfg of bullet_controller_one is
   for rtl
   end for;
end bullet_controller_one_rtl_cfg;
