configuration map_pass_controller_rtl_cfg of map_pass_controller is
   for rtl
   end for;
end map_pass_controller_rtl_cfg;
