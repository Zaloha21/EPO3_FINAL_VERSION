configuration bullet_pass_controller_rtl_cfg of bullet_pass_controller is
   for rtl
   end for;
end bullet_pass_controller_rtl_cfg;
