configuration map_switch_controller_rtl_cfg of map_switch_controller is
   for rtl
   end for;
end map_switch_controller_rtl_cfg;
