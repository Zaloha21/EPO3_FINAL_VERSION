configuration bullet_address_controller_rtl_cfg of bullet_address_controller is
   for rtl
   end for;
end bullet_address_controller_rtl_cfg;
