configuration bullet_pixel_mux_rtl_cfg of bullet_pixel_mux is
   for rtl
   end for;
end bullet_pixel_mux_rtl_cfg;
