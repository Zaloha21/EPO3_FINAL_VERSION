configuration pixel_mux_map_rtl_cfg of pixel_mux_map is
   for rtl
   end for;
end pixel_mux_map_rtl_cfg;
