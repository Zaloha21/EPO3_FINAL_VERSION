configuration vga_rgb_splitter_rtl_cfg of vga_rgb_splitter is
   for rtl
   end for;
end vga_rgb_splitter_rtl_cfg;
