configuration player_address_controller_rtl_cfg of player_address_controller is
   for rtl
   end for;
end player_address_controller_rtl_cfg;
