configuration rgb_rom_map_rtl_cfg of rgb_rom_map is
   for rtl
   end for;
end rgb_rom_map_rtl_cfg;
