configuration bullet_one_rgb_rom_rtl_cfg of bullet_one_rgb_rom is
   for rtl
   end for;
end bullet_one_rgb_rom_rtl_cfg;
