configuration bullet_two_rgb_rom_rtl_cfg of bullet_two_rgb_rom is
   for rtl
   end for;
end bullet_two_rgb_rom_rtl_cfg;
