configuration layer_mux_rtl_cfg of layer_mux is
   for rtl
   end for;
end layer_mux_rtl_cfg;
