configuration game_state_controller_rtl_cfg of game_state_controller is
   for rtl
   end for;
end game_state_controller_rtl_cfg;
