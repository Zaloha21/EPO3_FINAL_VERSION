configuration coordregister_behaviour_cfg of coordregister is
   for behaviour
   end for;
end coordregister_behaviour_cfg;
