configuration player_switch_controller_rtl_cfg of player_switch_controller is
   for rtl
   end for;
end player_switch_controller_rtl_cfg;
