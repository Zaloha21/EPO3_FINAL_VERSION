configuration pass_gate_rtl_cfg of pass_gate is
   for rtl
   end for;
end pass_gate_rtl_cfg;
