configuration player_pass_controller_rtl_cfg of player_pass_controller is
   for rtl
   end for;
end player_pass_controller_rtl_cfg;
