configuration player_one_rgb_rom_rtl_cfg of player_one_rgb_rom is
   for rtl
   end for;
end player_one_rgb_rom_rtl_cfg;
