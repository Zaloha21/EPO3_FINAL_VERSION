configuration rom_bus_rtl_cfg of rom_bus is
   for rtl
   end for;
end rom_bus_rtl_cfg;
