configuration vga_h_sync_gen_rtl_cfg of vga_h_sync_gen is
   for rtl
   end for;
end vga_h_sync_gen_rtl_cfg;
