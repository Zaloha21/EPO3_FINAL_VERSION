configuration map_pass_converter_rtl_cfg of map_pass_converter is
   for rtl
   end for;
end map_pass_converter_rtl_cfg;
