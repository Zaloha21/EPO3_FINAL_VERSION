configuration bullet_two_sprite_rom_rtl_cfg of bullet_two_sprite_rom is
   for rtl
   end for;
end bullet_two_sprite_rom_rtl_cfg;
