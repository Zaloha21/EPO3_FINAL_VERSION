configuration vga_v_sync_gen_rtl_cfg of vga_v_sync_gen is
   for rtl
   end for;
end vga_v_sync_gen_rtl_cfg;
