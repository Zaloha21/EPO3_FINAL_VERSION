configuration jumpregister_behaviour_cfg of jumpregister is
   for behaviour
   end for;
end jumpregister_behaviour_cfg;
