library IEEE;
use IEEE.std_logic_1164.all;

entity mes_chip_tb is
end entity mes_chip_tb;