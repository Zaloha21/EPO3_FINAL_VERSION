configuration bullet_controller_two_rtl_cfg of bullet_controller_two is
   for rtl
   end for;
end bullet_controller_two_rtl_cfg;
