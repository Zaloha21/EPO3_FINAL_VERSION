configuration map_address_controller_rtl_cfg of map_address_controller is
   for rtl
   end for;
end map_address_controller_rtl_cfg;
