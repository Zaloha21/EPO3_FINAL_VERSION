configuration map_rom_rtl_cfg of map_rom is
   for rtl
   end for;
end map_rom_rtl_cfg;
