configuration buttonreg_behaviour_cfg of buttonreg is
   for behaviour
   end for;
end buttonreg_behaviour_cfg;
