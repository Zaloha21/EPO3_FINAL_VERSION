configuration pixel_counter_rtl_cfg of pixel_counter is
   for rtl
   end for;
end pixel_counter_rtl_cfg;
