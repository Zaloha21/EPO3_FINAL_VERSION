configuration bullet_switch_controller_rtl_cfg of bullet_switch_controller is
   for rtl
   end for;
end bullet_switch_controller_rtl_cfg;
