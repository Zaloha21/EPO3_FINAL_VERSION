configuration dirregister_behaviour_cfg of dirregister is
   for behaviour
   end for;
end dirregister_behaviour_cfg;
